`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer:  Ndricim Rrapi & Argert Boja
// 
// Module Name:    SegmentDisplay
//
// Description: This module takes as inputs the current states of the elevators and the current state 
/*              of the person requesting the elevator. According to this data this module is implemented 
                in such a way that it will display these states in digits on Basys3 7Segment Display.
*/
// Project Name: Twin Elevator
//
// LED positions inside 7-segment
//    A 
//  F   B
//    G
//  E   C
//    D      DP

// digit positions on Basys3 :
// in3(left), in2, in1, in0(right)


module SegmentDisplay( input logic clk,input logic [3:0] csWire,csWire2,des1, des2,       // 4 values for 4 digits (decimal value)
                       output logic a, b, c, d, e, f, g, dp, //individual LED output for the 7-segment along with the digital point
                       output logic [3:0] an   // anode: 4-bit enable signal (active low)
                      );
 
    logic [3:0] in0, in1, in2,in3;
 
    // divide system clock (100Mhz for Basys3) by 2^N using a counter, which allows us to multiplex at lower speed
    localparam N = 18;
    logic [N-1:0] count = {N{1'b0}}; //initial value
    always@ (posedge clk)
        count <= count + 1;
    
     
    logic [3:0]digit_val; // 7-bit register to hold the current data on output
    logic [3:0]digit_en;  //register for enable vector
     
    always @*
    begin
        case (csWire)
            4'b0001: in0 <= csWire;
            4'b0010: in0 <= csWire;
            4'b0100: in0 <= 4'b0011;
            4'b1000: in0 <= 4'b0100;
            4'b0000 : in0 <= 4'b1001;
            default : in0 <= 4'b0000;
        endcase
       
         case (csWire2)
             4'b0001: in1 <= csWire2;
             4'b0010: in1 <= csWire2;
             4'b0100: in1 <= 4'b0011;
             4'b1000: in1 <= 4'b0100;
             4'b0000 : in1 <= 4'b1001;
             default:  in1 <= 4'b1000;
         endcase
                   
         case (des1)
              4'b0001: in2 <= des1;
              4'b0010: in2 <= des1;
              4'b0100: in2 <= 4'b0011;
              4'b1000: in2 <= 4'b0100;
              4'b0000 : in2 <= 4'b1001;
              default:  in2 <= 4'b1000;
         endcase
            
         case (des2)
               4'b0001: in3 <= des2;
               4'b0010: in3 <= des2;
               4'b0100: in3 <= 4'b0011;
               4'b1000: in3 <= 4'b0100;
               4'b0000 : in3 <= 4'b1001;
               default:  in3 <= 4'b1000;
          endcase
    end 
     
    always_comb
    begin
         digit_en = 4'b1111; //default
         digit_val = in0; //default
         
         case(count[N-1:N-2]) //using only the 2 MSB's of the counter 
            
           2'b00 :  //select first 7Seg.
            begin
             digit_val = in0;
             digit_en = 4'b1110;
            end
            
           2'b01:  //select second 7Seg.
            begin
             digit_val = in1;
             digit_en = 4'b1101;
            end
            
           2'b10:  //select third 7Seg.
            begin
             digit_val = in2;
             digit_en = 4'b1011;
            end
             
           2'b11:  //select forth 7Seg.
            begin
             digit_val = in3;
             digit_en = 4'b0111;
            end
         endcase
     end
     
    
    //Convert digit number to LED vector. LEDs are active low.
    logic [6:0] sseg_LEDs; 
    always_comb
     begin 
      sseg_LEDs = 7'b1111111; //default
      case(digit_val)
       4'd0 : sseg_LEDs = 7'b1000000; //to display 0
       4'd1 : sseg_LEDs = 7'b1111001; //to display 1
       4'd2 : sseg_LEDs = 7'b0100100; //to display 2
       4'd3 : sseg_LEDs = 7'b0110000; //to display 3
       4'd4 : sseg_LEDs = 7'b0011001; //to display 4
       4'd5 : sseg_LEDs = 7'b0010010; //to display 5
       4'd6 : sseg_LEDs = 7'b0000010; //to display 6
       4'd7 : sseg_LEDs = 7'b1111000; //to display 7
       4'd8 : sseg_LEDs = 7'b0000000; //to display 8
       4'd9 : sseg_LEDs = 7'b0010000; //to display 9
       default : sseg_LEDs = 7'b0111111; //dash
      endcase
     end
     
    assign an = digit_en; 
    assign {g, f, e, d, c, b, a} = sseg_LEDs; 
    assign dp = 1'b1; //turn dp off
     
endmodule
